module CNN(
    input wire clk,
    input wire rstn,
    input wire signed [31:0] din,
    output wire [9:0] classes,
    output wire done,  
);
endmodule