module conv_mix_tb ();
parameter cycle = 20;
reg clk;
reg rstn;
reg start_conv;
reg signed[31:0] image_in;
reg start_window;
reg state;
wire [159:0] taps;
reg weight_en;
reg weight_c;
wire [31:0] conv_result;
wire conv_done;
wire conv_ovalid;

integer fp_i;
integer count_w;

reg [10:0] cnt_line;
reg [10:0] cnt_conv;
reg signed [31:0] conv_result_r [0:599];

conv_mix conv_mix_inst(
    .clk(clk),
    .rstn(rstn),
    .start(start_conv),
    .weight_en(weight_en),
    .weight(weight_c),
    .din(image_in),
    .state(state),
    .ovalid(conv_ovalid),
    .done(conv_done),
    .dout(conv_result)
);

initial begin
    clk = 0;
    rstn = 0;
    state = 0;
    cnt_conv = 0;
    #20;
    rstn = 1;
    start_conv = 1;
    weight_en = 1;
    weight_c = 0;
end

initial begin
    fp_i = $fopen("/home/curry/code/curry_code_summay/rtl_works/BNN_on_fpga/test_image_txt.txt", "r");
end

always @(posedge clk) begin
    if(start_window == 1)
    begin
        count_w <= $fscanf(fp_i,"%b",image_in);
        cnt_line <= cnt_line + 1;
        if(cnt_line == 784) $display("image read done");
    end
end
integer i;
integer display_line = 0;
always @(posedge clk) begin
    if(conv_ovalid&& !conv_done)
    begin
        conv_result_r[cnt_conv] =  conv_result; 
        cnt_conv = cnt_conv + 1;
    end
    else begin
        if(conv_done) // 以24x24二维矩阵形式打印卷积结果
        begin
            conv_result_r[cnt_conv] =  conv_result; // 最后一个结果，conv_ovalid 和 conv_done均为 1
            //$display("cnt_conv: %d  ", cnt_conv);
            $display("conv complete");
            if(state == 0)
            begin
                for(i=0;i<576;i=i+1)
                begin 
                    if(i == 0) $write("%d :", display_line);
                    
                    $write("%d ", conv_result_r[i]); // $write 不会自动换行
                    
                    if((i+1)%24 == 0)// 添加行号并换行
                    begin
                        $display(" "); // 每行 24 个数据
                        display_line = display_line + 1;
                        $write("%d :", display_line);
                    end
                end	
            end
            else if(state == 1)
            begin
                for(i=0;i<64;i=i+1)
                begin
                    $display("%d", conv_result_r[i]);
                end	
            end
            
        end
    end
end

endmodule