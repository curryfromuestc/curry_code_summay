module window (
    input wire clk,
    input wire start,
    input wire [7:0] din,
    input wire state,
    output wire [39:0]taps
);

// 声明一个ram
reg [7:0] mem [139:0];

    
endmodule