module conv (
    ports
);
    
endmodule